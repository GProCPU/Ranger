`timescale  1ns/1ps

`include rv32.sv
`include ranger.sv


module control (
        input  logic clk,
        input  logic rst_n,
    );

endmodule
